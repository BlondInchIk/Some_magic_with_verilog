`timescale 1ns / 1ps
module SISO(input clk,b,output q);
wire w1,w2,w3;

d_ff dut1(
    .clk(clk),
    .d(b),
    .q(w1),
    .rst()
    );

d_ff dut2(
    .clk(clk),
    .d(w1),
    .q(w2),
    .rst()
    );
    
d_ff dut3(
    .clk(clk),
    .d(w2),
    .q(w3),
    .rst()
    );

d_ff dut4(
    .clk(clk),
    .d(w3),
    .q(q),
    .rst()
    );

endmodule

// d flip flop
module d_ff (
    input clk,    
    input d,      
    input rst,    
    output reg q);

    always @(posedge clk) 
    begin
    if (rst)
        q <= 1'b0;
    else
        q <= d;
    end

endmodule